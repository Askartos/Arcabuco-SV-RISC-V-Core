package arcabuco_system_config;
  parameter int NPADS=2;
endpackage
